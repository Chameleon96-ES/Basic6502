// CV96_QSYS.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module CV96_QSYS (
		output wire        hps_0_h2f_user0_clock_clk,      // hps_0_h2f_user0_clock.clk
		output wire        hps_0_h2f_user1_clock_clk,      // hps_0_h2f_user1_clock.clk
		input  wire        hps_io_hps_io_uart0_inst_RX,    //                hps_io.hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,    //                      .hps_io_uart0_inst_TX
		input  wire        hps_io_hps_io_uart0_inst_CTS,   //                      .hps_io_uart0_inst_CTS
		output wire        hps_io_hps_io_uart0_inst_RTS,   //                      .hps_io_uart0_inst_RTS
		inout  wire        hps_io_hps_io_gpio_inst_GPIO00, //                      .hps_io_gpio_inst_GPIO00
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09, //                      .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO14, //                      .hps_io_gpio_inst_GPIO14
		inout  wire        hps_io_hps_io_gpio_inst_GPIO15, //                      .hps_io_gpio_inst_GPIO15
		inout  wire        hps_io_hps_io_gpio_inst_GPIO16, //                      .hps_io_gpio_inst_GPIO16
		inout  wire        hps_io_hps_io_gpio_inst_GPIO17, //                      .hps_io_gpio_inst_GPIO17
		inout  wire        hps_io_hps_io_gpio_inst_GPIO18, //                      .hps_io_gpio_inst_GPIO18
		inout  wire        hps_io_hps_io_gpio_inst_GPIO19, //                      .hps_io_gpio_inst_GPIO19
		inout  wire        hps_io_hps_io_gpio_inst_GPIO22, //                      .hps_io_gpio_inst_GPIO22
		inout  wire        hps_io_hps_io_gpio_inst_GPIO23, //                      .hps_io_gpio_inst_GPIO23
		inout  wire        hps_io_hps_io_gpio_inst_GPIO24, //                      .hps_io_gpio_inst_GPIO24
		inout  wire        hps_io_hps_io_gpio_inst_GPIO25, //                      .hps_io_gpio_inst_GPIO25
		inout  wire        hps_io_hps_io_gpio_inst_GPIO26, //                      .hps_io_gpio_inst_GPIO26
		inout  wire        hps_io_hps_io_gpio_inst_GPIO27, //                      .hps_io_gpio_inst_GPIO27
		inout  wire        hps_io_hps_io_gpio_inst_GPIO28, //                      .hps_io_gpio_inst_GPIO28
		inout  wire        hps_io_hps_io_gpio_inst_GPIO29, //                      .hps_io_gpio_inst_GPIO29
		inout  wire        hps_io_hps_io_gpio_inst_GPIO30, //                      .hps_io_gpio_inst_GPIO30
		inout  wire        hps_io_hps_io_gpio_inst_GPIO31, //                      .hps_io_gpio_inst_GPIO31
		inout  wire        hps_io_hps_io_gpio_inst_GPIO32, //                      .hps_io_gpio_inst_GPIO32
		inout  wire        hps_io_hps_io_gpio_inst_GPIO33, //                      .hps_io_gpio_inst_GPIO33
		inout  wire        hps_io_hps_io_gpio_inst_GPIO34, //                      .hps_io_gpio_inst_GPIO34
		inout  wire        hps_io_hps_io_gpio_inst_GPIO37, //                      .hps_io_gpio_inst_GPIO37
		inout  wire        hps_io_hps_io_gpio_inst_GPIO44, //                      .hps_io_gpio_inst_GPIO44
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48, //                      .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53, //                      .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54, //                      .hps_io_gpio_inst_GPIO54
		output wire [13:0] memory_mem_a,                   //                memory.mem_a
		output wire [2:0]  memory_mem_ba,                  //                      .mem_ba
		output wire        memory_mem_ck,                  //                      .mem_ck
		output wire        memory_mem_ck_n,                //                      .mem_ck_n
		output wire        memory_mem_cke,                 //                      .mem_cke
		output wire        memory_mem_cs_n,                //                      .mem_cs_n
		output wire        memory_mem_ras_n,               //                      .mem_ras_n
		output wire        memory_mem_cas_n,               //                      .mem_cas_n
		output wire        memory_mem_we_n,                //                      .mem_we_n
		output wire        memory_mem_reset_n,             //                      .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                  //                      .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                 //                      .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,               //                      .mem_dqs_n
		output wire        memory_mem_odt,                 //                      .mem_odt
		output wire [1:0]  memory_mem_dm,                  //                      .mem_dm
		input  wire        memory_oct_rzqin                //                      .oct_rzqin
	);

	CV96_QSYS_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_user0_clk           (hps_0_h2f_user0_clock_clk),      // h2f_user0_clock.clk
		.h2f_user1_clk           (hps_0_h2f_user1_clock_clk),      // h2f_user1_clock.clk
		.mem_a                   (memory_mem_a),                   //          memory.mem_a
		.mem_ba                  (memory_mem_ba),                  //                .mem_ba
		.mem_ck                  (memory_mem_ck),                  //                .mem_ck
		.mem_ck_n                (memory_mem_ck_n),                //                .mem_ck_n
		.mem_cke                 (memory_mem_cke),                 //                .mem_cke
		.mem_cs_n                (memory_mem_cs_n),                //                .mem_cs_n
		.mem_ras_n               (memory_mem_ras_n),               //                .mem_ras_n
		.mem_cas_n               (memory_mem_cas_n),               //                .mem_cas_n
		.mem_we_n                (memory_mem_we_n),                //                .mem_we_n
		.mem_reset_n             (memory_mem_reset_n),             //                .mem_reset_n
		.mem_dq                  (memory_mem_dq),                  //                .mem_dq
		.mem_dqs                 (memory_mem_dqs),                 //                .mem_dqs
		.mem_dqs_n               (memory_mem_dqs_n),               //                .mem_dqs_n
		.mem_odt                 (memory_mem_odt),                 //                .mem_odt
		.mem_dm                  (memory_mem_dm),                  //                .mem_dm
		.oct_rzqin               (memory_oct_rzqin),               //                .oct_rzqin
		.hps_io_uart0_inst_RX    (hps_io_hps_io_uart0_inst_RX),    //          hps_io.hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX    (hps_io_hps_io_uart0_inst_TX),    //                .hps_io_uart0_inst_TX
		.hps_io_uart0_inst_CTS   (hps_io_hps_io_uart0_inst_CTS),   //                .hps_io_uart0_inst_CTS
		.hps_io_uart0_inst_RTS   (hps_io_hps_io_uart0_inst_RTS),   //                .hps_io_uart0_inst_RTS
		.hps_io_gpio_inst_GPIO00 (hps_io_hps_io_gpio_inst_GPIO00), //                .hps_io_gpio_inst_GPIO00
		.hps_io_gpio_inst_GPIO09 (hps_io_hps_io_gpio_inst_GPIO09), //                .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO14 (hps_io_hps_io_gpio_inst_GPIO14), //                .hps_io_gpio_inst_GPIO14
		.hps_io_gpio_inst_GPIO15 (hps_io_hps_io_gpio_inst_GPIO15), //                .hps_io_gpio_inst_GPIO15
		.hps_io_gpio_inst_GPIO16 (hps_io_hps_io_gpio_inst_GPIO16), //                .hps_io_gpio_inst_GPIO16
		.hps_io_gpio_inst_GPIO17 (hps_io_hps_io_gpio_inst_GPIO17), //                .hps_io_gpio_inst_GPIO17
		.hps_io_gpio_inst_GPIO18 (hps_io_hps_io_gpio_inst_GPIO18), //                .hps_io_gpio_inst_GPIO18
		.hps_io_gpio_inst_GPIO19 (hps_io_hps_io_gpio_inst_GPIO19), //                .hps_io_gpio_inst_GPIO19
		.hps_io_gpio_inst_GPIO22 (hps_io_hps_io_gpio_inst_GPIO22), //                .hps_io_gpio_inst_GPIO22
		.hps_io_gpio_inst_GPIO23 (hps_io_hps_io_gpio_inst_GPIO23), //                .hps_io_gpio_inst_GPIO23
		.hps_io_gpio_inst_GPIO24 (hps_io_hps_io_gpio_inst_GPIO24), //                .hps_io_gpio_inst_GPIO24
		.hps_io_gpio_inst_GPIO25 (hps_io_hps_io_gpio_inst_GPIO25), //                .hps_io_gpio_inst_GPIO25
		.hps_io_gpio_inst_GPIO26 (hps_io_hps_io_gpio_inst_GPIO26), //                .hps_io_gpio_inst_GPIO26
		.hps_io_gpio_inst_GPIO27 (hps_io_hps_io_gpio_inst_GPIO27), //                .hps_io_gpio_inst_GPIO27
		.hps_io_gpio_inst_GPIO28 (hps_io_hps_io_gpio_inst_GPIO28), //                .hps_io_gpio_inst_GPIO28
		.hps_io_gpio_inst_GPIO29 (hps_io_hps_io_gpio_inst_GPIO29), //                .hps_io_gpio_inst_GPIO29
		.hps_io_gpio_inst_GPIO30 (hps_io_hps_io_gpio_inst_GPIO30), //                .hps_io_gpio_inst_GPIO30
		.hps_io_gpio_inst_GPIO31 (hps_io_hps_io_gpio_inst_GPIO31), //                .hps_io_gpio_inst_GPIO31
		.hps_io_gpio_inst_GPIO32 (hps_io_hps_io_gpio_inst_GPIO32), //                .hps_io_gpio_inst_GPIO32
		.hps_io_gpio_inst_GPIO33 (hps_io_hps_io_gpio_inst_GPIO33), //                .hps_io_gpio_inst_GPIO33
		.hps_io_gpio_inst_GPIO34 (hps_io_hps_io_gpio_inst_GPIO34), //                .hps_io_gpio_inst_GPIO34
		.hps_io_gpio_inst_GPIO37 (hps_io_hps_io_gpio_inst_GPIO37), //                .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO44 (hps_io_hps_io_gpio_inst_GPIO44), //                .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48 (hps_io_hps_io_gpio_inst_GPIO48), //                .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53 (hps_io_hps_io_gpio_inst_GPIO53), //                .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54 (hps_io_hps_io_gpio_inst_GPIO54), //                .hps_io_gpio_inst_GPIO54
		.h2f_rst_n               ()                                //       h2f_reset.reset_n
	);

endmodule
